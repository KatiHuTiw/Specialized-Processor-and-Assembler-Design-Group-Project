module decoderModule()(
    input[8:0] binaryCode;
    output[4:0] opcode;
    output[1:0] operand1;
    output[1:0] operand2;
);