// program counter
// supports both relative and absolute jumps
// use either or both, as desired
module PC #(parameter D=12)(
  input reset,					// synchronous reset
        clk,
		  stall,
		  jump_en,             // jump enable (only relative)
  input       [D-1:0] target,	// how far/where to jump
  output logic[D-1:0] prog_ctr
);

  always_ff @(posedge clk)
    if(reset)
	  prog_ctr <= '0;
	else if(jump_en)
	  prog_ctr <= prog_ctr + 12'b1 + target;
	else if(stall)
	  prog_ctr <= prog_ctr + '0;
	else
	  prog_ctr <= prog_ctr + 12'b1;

endmodule
